// Configuration macros for systolic array parameters
`ifndef SYSTOLIC_CONFIG_VH
`define SYSTOLIC_CONFIG_VH

`ifndef SYSTOLIC_FRAC_WIDTH
`define SYSTOLIC_FRAC_WIDTH 15
`endif

`define SYSTOLIC_INPUT_WIDTH  16
`define SYSTOLIC_RESULT_WIDTH 16
`define SYSTOLIC_ADDR_WIDTH   10

`endif
